// Verilog test fixture created from schematic X:\EC311Lab1\Lab1.sch - Fri Feb 20 16:39:59 2015

`timescale 1ns / 1ps

module Lab1_Lab1_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Lab1 UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
